`timescale 1ns/1ns
module Shifter( in, inShift, Signal, out  ) ;

	input[31:0]		in ;
	input[31:0]		inShift ;
	input[5:0]		Signal ;
	output[31:0]	out ;
	
	wire[4:0]		shift ;
	wire[31:0]		temp ;
	wire[31:0]		temp2 ;
	wire[31:0]		temp3 ;
	wire[31:0]		temp4 ;
	wire[31:0]		temp5 ;
	
	// parameter SLL = 6'b000000 ;  // 左移???
	assign shift = inShift[4:0] ;
	
	// assign temp = ( shift[0] == 1'b1 ) ? {in[30:0],1'b0} : in ;
	// shift 1 bit
	assign temp[31] = shift[0] ? in[30] : in[31] ;
	assign temp[30] = shift[0] ? in[29] : in[30] ;
	assign temp[29] = shift[0] ? in[28] : in[29] ;
	assign temp[28] = shift[0] ? in[27] : in[28] ;
	assign temp[27] = shift[0] ? in[26] : in[27] ;
	assign temp[26] = shift[0] ? in[25] : in[26] ;	
	assign temp[25] = shift[0] ? in[24] : in[25] ;
	assign temp[24] = shift[0] ? in[23] : in[24] ;
	assign temp[23] = shift[0] ? in[22] : in[23] ;
	assign temp[22] = shift[0] ? in[21] : in[22] ;
	assign temp[21] = shift[0] ? in[20] : in[21] ;
	assign temp[20] = shift[0] ? in[19] : in[20] ;
	assign temp[19] = shift[0] ? in[18] : in[19] ;
	assign temp[18] = shift[0] ? in[17] : in[18] ;
	assign temp[17] = shift[0] ? in[16] : in[17] ;
	assign temp[16] = shift[0] ? in[15] : in[16] ;
	assign temp[15] = shift[0] ? in[14] : in[15] ;
	assign temp[14] = shift[0] ? in[13] : in[14] ;
	assign temp[13] = shift[0] ? in[12] : in[13] ;
	assign temp[12] = shift[0] ? in[11] : in[12] ;	
	assign temp[11] = shift[0] ? in[10] : in[11] ;
	assign temp[10] = shift[0] ? in[9] : in[10] ;
	assign temp[9] = shift[0] ? in[8] : in[9] ;
	assign temp[8] = shift[0] ? in[7] : in[8] ;
	assign temp[7] = shift[0] ? in[6] : in[7] ;
	assign temp[6] = shift[0] ? in[5] : in[6] ;
	assign temp[5] = shift[0] ? in[4] : in[5] ;
	assign temp[4] = shift[0] ? in[3] : in[4] ;
	assign temp[3] = shift[0] ? in[2] : in[3] ;
	assign temp[2] = shift[0] ? in[1] : in[2] ;
	assign temp[1] = shift[0] ? in[0] : in[1] ;
	assign temp[0] = shift[0] ? 1'b0 : in[0] ;
	// assign temp2 = ( shift[1] == 1'b1 ) ? {temp[29:0],2'b0} : temp ;
	// shift 2 bit
	assign temp2[31] = shift[1] ? temp[29] : temp[31] ;
	assign temp2[30] = shift[1] ? temp[28] : temp[30] ;
	assign temp2[29] = shift[1] ? temp[27] : temp[29] ;
	assign temp2[28] = shift[1] ? temp[26] : temp[28] ;
	assign temp2[27] = shift[1] ? temp[25] : temp[27] ;
	assign temp2[26] = shift[1] ? temp[24] : temp[26] ;	
	assign temp2[25] = shift[1] ? temp[23] : temp[25] ;
	assign temp2[24] = shift[1] ? temp[22] : temp[24] ;
	assign temp2[23] = shift[1] ? temp[21] : temp[23] ;
	assign temp2[22] = shift[1] ? temp[20] : temp[22] ;
	assign temp2[21] = shift[1] ? temp[19] : temp[21] ;
	assign temp2[20] = shift[1] ? temp[18] : temp[20] ;
	assign temp2[19] = shift[1] ? temp[17] : temp[19] ;
	assign temp2[18] = shift[1] ? temp[16] : temp[18] ;
	assign temp2[17] = shift[1] ? temp[15] : temp[17] ;
	assign temp2[16] = shift[1] ? temp[14] : temp[16] ;
	assign temp2[15] = shift[1] ? temp[13] : temp[15] ;
	assign temp2[14] = shift[1] ? temp[12] : temp[14] ;
	assign temp2[13] = shift[1] ? temp[11] : temp[13] ;
	assign temp2[12] = shift[1] ? temp[10] : temp[12] ;	
	assign temp2[11] = shift[1] ? temp[9] : temp[11] ;
	assign temp2[10] = shift[1] ? temp[8] : temp[10] ;
	assign temp2[9] = shift[1] ? temp[7] : temp[9] ;
	assign temp2[8] = shift[1] ? temp[6] : temp[8] ;
	assign temp2[7] = shift[1] ? temp[5] : temp[7] ;
	assign temp2[6] = shift[1] ? temp[4] : temp[6] ;
	assign temp2[5] = shift[1] ? temp[3] : temp[5] ;
	assign temp2[4] = shift[1] ? temp[2] : temp[4] ;
	assign temp2[3] = shift[1] ? temp[1] : temp[3] ;
	assign temp2[2] = shift[1] ? temp[0] : temp[2] ;
	assign temp2[1] = shift[1] ? 1'b0 : temp[1] ;
	assign temp2[0] = shift[1] ? 1'b0 : temp[0] ;
	// assign temp3 = ( shift[2] == 1'b1 ) ? {temp2[27:0],4'b0} : temp2 ;
	// shift 4 bit
	assign temp3[31] = shift[2] ? temp2[27] : temp2[31] ;
	assign temp3[30] = shift[2] ? temp2[26] : temp2[30] ;
	assign temp3[29] = shift[2] ? temp2[25] : temp2[29] ;
	assign temp3[28] = shift[2] ? temp2[24] : temp2[28] ;
	assign temp3[27] = shift[2] ? temp2[23] : temp2[27] ;
	assign temp3[26] = shift[2] ? temp2[22] : temp2[26] ;	
	assign temp3[25] = shift[2] ? temp2[21] : temp2[25] ;
	assign temp3[24] = shift[2] ? temp2[20] : temp2[24] ;
	assign temp3[23] = shift[2] ? temp2[19] : temp2[23] ;
	assign temp3[22] = shift[2] ? temp2[18] : temp2[22] ;
	assign temp3[21] = shift[2] ? temp2[17] : temp2[21] ;
	assign temp3[20] = shift[2] ? temp2[16] : temp2[20] ;
	assign temp3[19] = shift[2] ? temp2[15] : temp2[19] ;
	assign temp3[18] = shift[2] ? temp2[14] : temp2[18] ;
	assign temp3[17] = shift[2] ? temp2[13] : temp2[17] ;
	assign temp3[16] = shift[2] ? temp2[12] : temp2[16] ;
	assign temp3[15] = shift[2] ? temp2[11] : temp2[15] ;
	assign temp3[14] = shift[2] ? temp2[10] : temp2[14] ;
	assign temp3[13] = shift[2] ? temp2[9] : temp2[13] ;
	assign temp3[12] = shift[2] ? temp2[8] : temp2[12] ;	
	assign temp3[11] = shift[2] ? temp2[7] : temp2[11] ;
	assign temp3[10] = shift[2] ? temp2[6] : temp2[10] ;
	assign temp3[9] = shift[2] ? temp2[5] : temp2[9] ;
	assign temp3[8] = shift[2] ? temp2[4] : temp2[8] ;
	assign temp3[7] = shift[2] ? temp2[3] : temp2[7] ;
	assign temp3[6] = shift[2] ? temp2[2] : temp2[6] ;
	assign temp3[5] = shift[2] ? temp2[1] : temp2[5] ;
	assign temp3[4] = shift[2] ? temp2[0] : temp2[4] ;
	assign temp3[3] = shift[2] ? 1'b0 : temp2[3] ;
	assign temp3[2] = shift[2] ? 1'b0 : temp2[2] ;
	assign temp3[1] = shift[2] ? 1'b0 : temp2[1] ;
	assign temp3[0] = shift[2] ? 1'b0 : temp2[0] ;
	// assign temp4 = ( shift[3] == 1'b1 ) ? {temp3[23:0],8'b0} : temp3 ;
	// shift 8 bit
	assign temp4[31] = shift[3] ? temp3[23] : temp3[31] ;
	assign temp4[30] = shift[3] ? temp3[22] : temp3[30] ;
	assign temp4[29] = shift[3] ? temp3[21] : temp3[29] ;
	assign temp4[28] = shift[3] ? temp3[20] : temp3[28] ;
	assign temp4[27] = shift[3] ? temp3[19] : temp3[27] ;
	assign temp4[26] = shift[3] ? temp3[18] : temp3[26] ;	
	assign temp4[25] = shift[3] ? temp3[17] : temp3[25] ;
	assign temp4[24] = shift[3] ? temp3[16] : temp3[24] ;
	assign temp4[23] = shift[3] ? temp3[15] : temp3[23] ;
	assign temp4[22] = shift[3] ? temp3[14] : temp3[22] ;
	assign temp4[21] = shift[3] ? temp3[13] : temp3[21] ;
	assign temp4[20] = shift[3] ? temp3[12] : temp3[20] ;
	assign temp4[19] = shift[3] ? temp3[11] : temp3[19] ;
	assign temp4[18] = shift[3] ? temp3[10] : temp3[18] ;
	assign temp4[17] = shift[3] ? temp3[9] : temp3[17] ;
	assign temp4[16] = shift[3] ? temp3[8] : temp3[16] ;
	assign temp4[15] = shift[3] ? temp3[7] : temp3[15] ;
	assign temp4[14] = shift[3] ? temp3[6] : temp3[14] ;
	assign temp4[13] = shift[3] ? temp3[5] : temp3[13] ;
	assign temp4[12] = shift[3] ? temp3[4] : temp3[12] ;	
	assign temp4[11] = shift[3] ? temp3[3] : temp3[11] ;
	assign temp4[10] = shift[3] ? temp3[2] : temp3[10] ;
	assign temp4[9] = shift[3] ? temp3[1] : temp3[9] ;
	assign temp4[8] = shift[3] ? temp3[0] : temp3[8] ;
	assign temp4[7] = shift[3] ? 1'b0 : temp3[7] ;
	assign temp4[6] = shift[3] ? 1'b0 : temp3[6] ;
	assign temp4[5] = shift[3] ? 1'b0 : temp3[5] ;
	assign temp4[4] = shift[3] ? 1'b0 : temp3[4] ;
	assign temp4[3] = shift[3] ? 1'b0 : temp3[3] ;
	assign temp4[2] = shift[3] ? 1'b0 : temp3[2] ;
	assign temp4[1] = shift[3] ? 1'b0 : temp3[1] ;
	assign temp4[0] = shift[3] ? 1'b0 : temp3[0] ;
	// assign temp5 = ( shift[4] == 1'b1 ) ? {temp4[15:0],16'b0} : temp4 ;
	// shift 16 bit
	assign temp5[31] = shift[4] ? temp4[15] : temp4[31] ;
	assign temp5[30] = shift[4] ? temp4[14] : temp4[30] ;
	assign temp5[29] = shift[4] ? temp4[13] : temp4[29] ;
	assign temp5[28] = shift[4] ? temp4[12] : temp4[28] ;
	assign temp5[27] = shift[4] ? temp4[11] : temp4[27] ;
	assign temp5[26] = shift[4] ? temp4[10] : temp4[26] ;	
	assign temp5[25] = shift[4] ? temp4[9] : temp4[25] ;
	assign temp5[24] = shift[4] ? temp4[8] : temp4[24] ;
	assign temp5[23] = shift[4] ? temp4[7] : temp4[23] ;
	assign temp5[22] = shift[4] ? temp4[6] : temp4[22] ;
	assign temp5[21] = shift[4] ? temp4[5] : temp4[21] ;
	assign temp5[20] = shift[4] ? temp4[4] : temp4[20] ;
	assign temp5[19] = shift[4] ? temp4[3] : temp4[19] ;
	assign temp5[18] = shift[4] ? temp4[2] : temp4[18] ;
	assign temp5[17] = shift[4] ? temp4[1] : temp4[17] ;
	assign temp5[16] = shift[4] ? temp4[0] : temp4[16] ;
	assign temp5[15] = shift[4] ? 1'b0 : temp4[15] ;
	assign temp5[14] = shift[4] ? 1'b0 : temp4[14] ;
	assign temp5[13] = shift[4] ? 1'b0 : temp4[13] ;
	assign temp5[12] = shift[4] ? 1'b0 : temp4[12] ;	
	assign temp5[11] = shift[4] ? 1'b0 : temp4[11] ;
	assign temp5[10] = shift[4] ? 1'b0 : temp4[10] ;
	assign temp5[9] = shift[4] ? 1'b0 : temp4[9] ;
	assign temp5[8] = shift[4] ? 1'b0 : temp4[8] ;
	assign temp5[7] = shift[4] ? 1'b0 : temp4[7] ;
	assign temp5[6] = shift[4] ? 1'b0 : temp4[6] ;
	assign temp5[5] = shift[4] ? 1'b0 : temp4[5] ;
	assign temp5[4] = shift[4] ? 1'b0 : temp4[4] ;
	assign temp5[3] = shift[4] ? 1'b0 : temp4[3] ;
	assign temp5[2] = shift[4] ? 1'b0 : temp4[2] ;
	assign temp5[1] = shift[4] ? 1'b0 : temp4[1] ;
	assign temp5[0] = shift[4] ? 1'b0 : temp4[0] ;
	
	assign out = ( Signal == 6'b000000 ) ? (( inShift > 31 ) ? 32'b0 : temp5 ) : out ;

	
endmodule